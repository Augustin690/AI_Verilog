`include "nn_layers.sv"

module simple_nn_top#(
    parameter N_INPUTS = 100,
    parameter N_LAYER1 = 32,
    parameter N_LAYER2 = 16,
    parameter N_LAYER3 = 10
)(
    input logic signed [15:0] input_vec [N_INPUTS],
    output logic [$clog2(N_LAYER3)-1:0] prediction
);
    // Placeholder weights (to be filled with real values)
    logic signed [15:0] weights1 [100][32];
    initial begin 
        weights1[0] = '{16'sd131, 16'sd88, 16'sd49, 16'sd86, -16'sd118, 16'sd61, 16'sd117, 16'sd71, -16'sd56, 16'sd11, 16'sd29, -16'sd50, 16'sd22, 16'sd110, 16'sd57, 16'sd16, 16'sd73, 16'sd70, 16'sd13, -16'sd127, 16'sd106, -16'sd1, -16'sd16, 16'sd91, 16'sd92, -16'sd79, -16'sd67, -16'sd95, 16'sd101, -16'sd43, -16'sd151, 16'sd88};
        weights1[1] = '{16'sd126, 16'sd22, -16'sd50, 16'sd6, -16'sd68, 16'sd40, 16'sd34, 16'sd24, -16'sd23, 16'sd41, -16'sd9, -16'sd47, 16'sd109, 16'sd45, 16'sd89, -16'sd7, -16'sd3, 16'sd114, 16'sd2, -16'sd118, 16'sd72, 16'sd16, -16'sd66, 16'sd158, 16'sd42, -16'sd99, -16'sd28, -16'sd34, 16'sd155, -16'sd67, -16'sd100, 16'sd56};
        weights1[2] = '{16'sd32, -16'sd43, -16'sd71, -16'sd27, -16'sd65, -16'sd24, 16'sd145, -16'sd25, -16'sd104, 16'sd49, 16'sd87, 16'sd51, 16'sd48, -16'sd28, -16'sd59, 16'sd153, -16'sd88, 16'sd6, -16'sd6, -16'sd106, 16'sd131, -16'sd89, -16'sd110, 16'sd32, 16'sd69, 16'sd30, 16'sd49, 16'sd41, 16'sd212, -16'sd15, -16'sd70, 16'sd56};
        weights1[3] = '{16'sd119, -16'sd182, 16'sd78, -16'sd158, 16'sd13, -16'sd11, 16'sd138, 16'sd120, 16'sd27, 16'sd131, 16'sd31, 16'sd108, -16'sd105, 16'sd118, 16'sd2, 16'sd188, -16'sd88, -16'sd182, -16'sd205, -16'sd134, 16'sd141, 16'sd146, -16'sd110, -16'sd65, 16'sd35, 16'sd123, 16'sd157, 16'sd59, 16'sd188, 16'sd45, -16'sd9, -16'sd124};
        weights1[4] = '{16'sd39, -16'sd168, 16'sd34, -16'sd199, -16'sd53, -16'sd107, 16'sd115, 16'sd88, 16'sd91, 16'sd18, 16'sd47, 16'sd79, -16'sd77, -16'sd27, -16'sd177, 16'sd118, -16'sd126, -16'sd98, -16'sd140, -16'sd200, 16'sd95, 16'sd99, -16'sd109, -16'sd57, 16'sd78, 16'sd131, 16'sd213, 16'sd30, 16'sd92, 16'sd112, -16'sd104, -16'sd183};
        weights1[5] = '{16'sd81, -16'sd156, 16'sd89, -16'sd106, 16'sd19, -16'sd176, 16'sd62, 16'sd53, 16'sd102, 16'sd9, 16'sd43, 16'sd81, -16'sd104, 16'sd33, -16'sd72, 16'sd100, 16'sd28, -16'sd50, -16'sd76, -16'sd140, -16'sd10, 16'sd24, -16'sd144, -16'sd49, 16'sd20, 16'sd89, 16'sd147, 16'sd25, 16'sd41, 16'sd26, -16'sd152, -16'sd102};
        weights1[6] = '{16'sd12, -16'sd91, 16'sd129, -16'sd170, 16'sd52, -16'sd61, 16'sd106, 16'sd62, -16'sd18, -16'sd11, -16'sd53, 16'sd27, -16'sd93, 16'sd128, 16'sd24, 16'sd98, -16'sd75, 16'sd117, -16'sd66, -16'sd63, 16'sd100, 16'sd75, -16'sd170, -16'sd54, 16'sd2, 16'sd89, 16'sd157, 16'sd110, 16'sd33, 16'sd118, -16'sd56, -16'sd69};
        weights1[7] = '{16'sd101, -16'sd186, 16'sd107, -16'sd109, 16'sd126, 16'sd12, 16'sd67, 16'sd101, -16'sd16, 16'sd17, -16'sd82, -16'sd46, -16'sd109, 16'sd146, 16'sd135, 16'sd159, -16'sd46, 16'sd74, -16'sd146, -16'sd50, 16'sd129, 16'sd110, -16'sd121, 16'sd21, -16'sd184, 16'sd61, 16'sd134, 16'sd148, 16'sd106, 16'sd204, -16'sd35, -16'sd158};
        weights1[8] = '{16'sd92, -16'sd83, 16'sd122, -16'sd58, 16'sd82, 16'sd34, 16'sd99, 16'sd24, -16'sd9, 16'sd56, -16'sd138, -16'sd92, -16'sd108, 16'sd167, 16'sd153, 16'sd152, -16'sd20, 16'sd18, -16'sd76, 16'sd121, 16'sd86, 16'sd146, -16'sd102, -16'sd22, -16'sd176, 16'sd13, 16'sd92, 16'sd103, 16'sd59, 16'sd146, 16'sd66, -16'sd169};
        weights1[9] = '{-16'sd167, -16'sd72, -16'sd180, -16'sd38, 16'sd61, 16'sd145, 16'sd89, -16'sd93, 16'sd129, -16'sd127, -16'sd107, 16'sd70, -16'sd99, 16'sd146, 16'sd114, 16'sd49, 16'sd132, -16'sd48, 16'sd154, 16'sd165, -16'sd78, 16'sd122, -16'sd76, -16'sd148, -16'sd129, 16'sd102, -16'sd98, 16'sd133, 16'sd107, 16'sd39, -16'sd19, -16'sd182};
        weights1[10] = '{16'sd79, 16'sd103, 16'sd2, 16'sd0, -16'sd87, 16'sd49, 16'sd109, 16'sd118, -16'sd82, 16'sd8, 16'sd85, -16'sd21, 16'sd111, 16'sd97, 16'sd118, 16'sd16, 16'sd99, 16'sd70, 16'sd64, -16'sd194, 16'sd27, 16'sd0, -16'sd4, 16'sd137, 16'sd74, -16'sd127, -16'sd129, -16'sd114, 16'sd91, -16'sd31, -16'sd142, 16'sd31};
        weights1[11] = '{16'sd117, 16'sd8, -16'sd2, 16'sd58, -16'sd51, -16'sd13, 16'sd74, 16'sd116, -16'sd64, -16'sd61, -16'sd16, -16'sd28, 16'sd44, -16'sd12, 16'sd95, 16'sd72, 16'sd76, 16'sd88, 16'sd80, -16'sd118, -16'sd42, -16'sd35, -16'sd7, 16'sd101, 16'sd123, -16'sd153, -16'sd55, -16'sd197, 16'sd151, -16'sd29, -16'sd159, 16'sd77};
        weights1[12] = '{16'sd33, -16'sd42, 16'sd22, -16'sd48, -16'sd11, -16'sd142, 16'sd122, 16'sd12, -16'sd80, 16'sd32, 16'sd45, 16'sd100, 16'sd130, -16'sd44, 16'sd13, 16'sd70, 16'sd40, 16'sd102, 16'sd54, -16'sd69, -16'sd18, -16'sd74, -16'sd83, 16'sd63, 16'sd38, -16'sd53, 16'sd17, -16'sd54, 16'sd105, 16'sd23, -16'sd96, 16'sd92};
        weights1[13] = '{16'sd82, -16'sd21, -16'sd18, 16'sd7, -16'sd27, -16'sd161, 16'sd69, 16'sd27, -16'sd24, 16'sd45, 16'sd3, 16'sd54, 16'sd94, 16'sd25, -16'sd69, 16'sd19, -16'sd54, 16'sd6, 16'sd58, -16'sd27, -16'sd20, -16'sd94, -16'sd80, 16'sd34, 16'sd33, 16'sd83, -16'sd51, 16'sd4, 16'sd124, -16'sd40, -16'sd12, 16'sd104};
        weights1[14] = '{16'sd73, 16'sd19, 16'sd20, -16'sd36, 16'sd40, -16'sd88, 16'sd53, 16'sd0, 16'sd22, 16'sd19, 16'sd74, 16'sd12, 16'sd68, -16'sd142, -16'sd41, -16'sd9, 16'sd8, -16'sd172, 16'sd81, -16'sd6, -16'sd3, -16'sd68, -16'sd91, 16'sd56, -16'sd11, 16'sd58, -16'sd82, 16'sd27, 16'sd40, -16'sd19, 16'sd11, 16'sd157};
        weights1[15] = '{16'sd59, 16'sd35, 16'sd70, -16'sd79, 16'sd48, -16'sd28, 16'sd24, 16'sd11, 16'sd147, 16'sd13, 16'sd54, 16'sd76, 16'sd45, -16'sd36, 16'sd121, 16'sd45, 16'sd81, -16'sd121, 16'sd49, 16'sd58, -16'sd31, -16'sd30, -16'sd91, 16'sd16, 16'sd48, 16'sd53, -16'sd14, -16'sd5, 16'sd30, -16'sd62, -16'sd75, -16'sd6};
        weights1[16] = '{16'sd50, -16'sd54, 16'sd90, -16'sd44, 16'sd108, -16'sd53, 16'sd48, -16'sd7, 16'sd70, 16'sd4, -16'sd36, 16'sd100, 16'sd21, 16'sd13, 16'sd68, -16'sd10, -16'sd16, -16'sd102, -16'sd4, 16'sd53, -16'sd56, 16'sd32, -16'sd64, 16'sd1, 16'sd10, 16'sd54, -16'sd28, 16'sd91, 16'sd91, 16'sd3, -16'sd44, -16'sd47};
        weights1[17] = '{16'sd6, -16'sd113, 16'sd78, -16'sd35, 16'sd63, -16'sd81, 16'sd67, -16'sd29, 16'sd66, -16'sd87, -16'sd30, 16'sd50, -16'sd69, 16'sd22, 16'sd62, 16'sd112, 16'sd28, -16'sd19, 16'sd61, 16'sd26, -16'sd38, 16'sd43, -16'sd63, -16'sd7, 16'sd14, 16'sd67, -16'sd1, 16'sd77, -16'sd1, 16'sd71, -16'sd49, -16'sd91};
        weights1[18] = '{-16'sd24, -16'sd141, 16'sd34, -16'sd103, 16'sd91, -16'sd60, -16'sd18, 16'sd39, 16'sd30, -16'sd1, -16'sd115, 16'sd14, -16'sd86, 16'sd131, 16'sd115, 16'sd124, 16'sd30, -16'sd101, 16'sd13, 16'sd41, -16'sd1, 16'sd44, -16'sd55, -16'sd67, -16'sd68, 16'sd36, 16'sd40, 16'sd68, 16'sd37, 16'sd98, -16'sd24, -16'sd156};
        weights1[19] = '{-16'sd26, -16'sd15, -16'sd121, -16'sd21, 16'sd87, 16'sd47, 16'sd100, -16'sd21, 16'sd113, -16'sd69, -16'sd96, 16'sd24, 16'sd38, 16'sd82, 16'sd94, 16'sd26, -16'sd35, -16'sd101, 16'sd110, 16'sd47, -16'sd80, 16'sd21, -16'sd73, -16'sd127, -16'sd119, 16'sd128, -16'sd34, 16'sd72, 16'sd9, 16'sd36, 16'sd44, -16'sd39};
        weights1[20] = '{16'sd101, 16'sd62, 16'sd17, 16'sd80, -16'sd73, 16'sd50, -16'sd16, 16'sd93, -16'sd118, 16'sd171, 16'sd108, -16'sd76, 16'sd61, 16'sd150, 16'sd88, 16'sd63, 16'sd63, 16'sd48, 16'sd48, -16'sd172, 16'sd157, 16'sd26, 16'sd63, 16'sd152, 16'sd55, -16'sd103, -16'sd119, -16'sd109, 16'sd106, -16'sd74, -16'sd104, -16'sd4};
        weights1[21] = '{16'sd143, 16'sd11, 16'sd83, 16'sd13, -16'sd92, -16'sd41, 16'sd47, 16'sd69, -16'sd37, -16'sd19, 16'sd61, -16'sd24, 16'sd118, 16'sd94, 16'sd34, 16'sd21, 16'sd51, 16'sd3, 16'sd46, -16'sd109, 16'sd6, 16'sd3, 16'sd25, 16'sd165, 16'sd30, -16'sd82, -16'sd53, -16'sd102, 16'sd139, -16'sd58, -16'sd170, 16'sd31};
        weights1[22] = '{16'sd95, 16'sd56, -16'sd46, -16'sd32, -16'sd28, -16'sd4, 16'sd87, 16'sd3, 16'sd36, 16'sd72, 16'sd49, -16'sd58, 16'sd12, 16'sd82, 16'sd121, 16'sd0, 16'sd71, 16'sd77, 16'sd27, -16'sd41, 16'sd57, -16'sd17, -16'sd3, 16'sd18, 16'sd6, -16'sd5, -16'sd122, -16'sd35, 16'sd138, 16'sd45, -16'sd49, 16'sd4};
        weights1[23] = '{16'sd64, 16'sd26, -16'sd61, 16'sd73, 16'sd13, 16'sd15, 16'sd27, -16'sd1, -16'sd18, 16'sd79, 16'sd41, -16'sd30, 16'sd114, 16'sd119, 16'sd81, 16'sd48, 16'sd65, 16'sd57, 16'sd38, 16'sd1, 16'sd127, 16'sd48, 16'sd21, 16'sd63, 16'sd25, 16'sd44, -16'sd144, -16'sd12, 16'sd23, 16'sd63, 16'sd39, 16'sd57};
        weights1[24] = '{16'sd4, 16'sd18, -16'sd25, 16'sd94, 16'sd2, 16'sd22, 16'sd30, -16'sd39, 16'sd37, 16'sd84, 16'sd59, 16'sd28, 16'sd97, 16'sd33, 16'sd22, 16'sd18, 16'sd48, -16'sd130, 16'sd99, 16'sd65, 16'sd3, 16'sd53, 16'sd83, 16'sd14, 16'sd37, -16'sd41, -16'sd72, 16'sd4, 16'sd13, 16'sd50, 16'sd54, 16'sd94};
        weights1[25] = '{16'sd96, 16'sd80, -16'sd24, 16'sd76, 16'sd127, -16'sd17, 16'sd110, -16'sd48, 16'sd21, 16'sd14, 16'sd62, 16'sd85, 16'sd52, 16'sd9, -16'sd26, 16'sd36, 16'sd40, -16'sd11, 16'sd80, 16'sd99, 16'sd44, -16'sd27, 16'sd118, 16'sd31, 16'sd9, -16'sd60, 16'sd18, 16'sd27, -16'sd87, -16'sd54, 16'sd141, 16'sd152};
        weights1[26] = '{16'sd68, 16'sd128, 16'sd80, 16'sd69, 16'sd59, 16'sd62, 16'sd8, 16'sd3, 16'sd84, -16'sd4, 16'sd89, 16'sd33, 16'sd53, 16'sd69, 16'sd77, -16'sd58, 16'sd73, 16'sd44, 16'sd27, 16'sd136, 16'sd39, 16'sd12, 16'sd10, 16'sd44, 16'sd37, 16'sd3, 16'sd52, 16'sd52, -16'sd18, -16'sd3, 16'sd102, 16'sd147};
        weights1[27] = '{16'sd0, 16'sd47, 16'sd128, -16'sd16, 16'sd52, 16'sd102, -16'sd35, -16'sd30, 16'sd64, 16'sd0, 16'sd100, 16'sd32, 16'sd40, 16'sd38, 16'sd114, 16'sd30, 16'sd63, 16'sd5, 16'sd58, 16'sd82, 16'sd3, 16'sd57, -16'sd11, 16'sd43, -16'sd3, -16'sd5, 16'sd2, 16'sd65, -16'sd8, 16'sd41, 16'sd78, -16'sd1};
        weights1[28] = '{-16'sd43, -16'sd23, 16'sd65, -16'sd66, 16'sd85, 16'sd73, -16'sd1, -16'sd80, 16'sd57, 16'sd36, -16'sd78, -16'sd23, -16'sd90, 16'sd83, 16'sd42, 16'sd83, 16'sd78, -16'sd20, -16'sd52, 16'sd39, 16'sd4, 16'sd116, -16'sd62, -16'sd28, -16'sd103, 16'sd54, -16'sd41, 16'sd93, 16'sd7, 16'sd15, 16'sd36, -16'sd58};
        weights1[29] = '{-16'sd65, -16'sd39, -16'sd123, -16'sd21, 16'sd113, 16'sd84, 16'sd192, 16'sd6, 16'sd121, -16'sd118, -16'sd83, 16'sd76, -16'sd126, 16'sd44, 16'sd77, 16'sd129, -16'sd8, -16'sd78, 16'sd106, 16'sd98, -16'sd62, 16'sd99, -16'sd31, -16'sd139, -16'sd81, 16'sd66, -16'sd28, 16'sd108, 16'sd40, 16'sd123, -16'sd28, -16'sd144};
        weights1[30] = '{16'sd59, 16'sd126, 16'sd115, -16'sd23, -16'sd130, -16'sd138, -16'sd11, 16'sd116, -16'sd39, 16'sd286, 16'sd217, -16'sd36, 16'sd167, 16'sd96, -16'sd25, -16'sd170, 16'sd185, -16'sd287, 16'sd66, -16'sd186, -16'sd22, -16'sd156, 16'sd70, 16'sd134, 16'sd214, -16'sd34, -16'sd113, -16'sd109, 16'sd73, -16'sd263, -16'sd155, 16'sd108};
        weights1[31] = '{16'sd16, 16'sd59, 16'sd77, -16'sd6, -16'sd122, -16'sd58, 16'sd58, 16'sd73, -16'sd61, 16'sd0, 16'sd73, 16'sd17, 16'sd63, 16'sd66, 16'sd105, -16'sd105, 16'sd15, -16'sd121, 16'sd49, -16'sd143, 16'sd57, -16'sd100, 16'sd35, 16'sd113, 16'sd35, -16'sd15, -16'sd164, -16'sd110, 16'sd161, -16'sd123, -16'sd110, -16'sd55};
        weights1[32] = '{16'sd44, 16'sd47, -16'sd20, 16'sd4, -16'sd95, -16'sd48, 16'sd55, -16'sd102, 16'sd63, 16'sd43, 16'sd64, -16'sd37, 16'sd81, 16'sd52, -16'sd1, 16'sd42, -16'sd2, 16'sd113, 16'sd84, -16'sd12, 16'sd82, -16'sd21, 16'sd21, 16'sd27, -16'sd2, 16'sd21, -16'sd197, -16'sd17, 16'sd72, 16'sd43, -16'sd13, -16'sd78};
        weights1[33] = '{-16'sd41, 16'sd75, -16'sd12, -16'sd14, -16'sd64, 16'sd25, 16'sd4, -16'sd117, 16'sd74, 16'sd100, 16'sd56, 16'sd26, 16'sd53, 16'sd110, 16'sd33, 16'sd25, -16'sd30, -16'sd80, 16'sd70, 16'sd62, 16'sd51, 16'sd54, 16'sd42, 16'sd115, -16'sd58, 16'sd58, -16'sd17, 16'sd57, -16'sd42, 16'sd84, 16'sd60, -16'sd93};
        weights1[34] = '{-16'sd40, 16'sd57, -16'sd128, 16'sd85, 16'sd50, 16'sd27, -16'sd42, -16'sd97, 16'sd0, 16'sd104, -16'sd34, 16'sd37, -16'sd80, -16'sd13, 16'sd15, 16'sd91, -16'sd5, -16'sd196, 16'sd85, 16'sd97, -16'sd17, 16'sd51, 16'sd119, 16'sd156, -16'sd49, 16'sd37, 16'sd73, 16'sd25, -16'sd7, -16'sd32, 16'sd98, -16'sd44};
        weights1[35] = '{-16'sd72, 16'sd103, -16'sd206, 16'sd98, 16'sd16, 16'sd67, -16'sd75, 16'sd102, 16'sd7, 16'sd26, 16'sd55, 16'sd27, -16'sd1, -16'sd49, 16'sd31, 16'sd19, 16'sd37, 16'sd92, -16'sd3, 16'sd17, 16'sd41, -16'sd49, 16'sd131, 16'sd90, 16'sd113, -16'sd54, -16'sd47, -16'sd62, 16'sd80, -16'sd197, -16'sd29, 16'sd58};
        weights1[36] = '{16'sd77, 16'sd67, 16'sd143, 16'sd74, -16'sd114, 16'sd126, 16'sd51, 16'sd45, 16'sd13, 16'sd116, -16'sd8, 16'sd0, -16'sd32, 16'sd39, 16'sd63, -16'sd121, 16'sd85, 16'sd170, -16'sd31, 16'sd31, 16'sd43, 16'sd23, 16'sd27, 16'sd74, 16'sd41, -16'sd12, -16'sd37, -16'sd92, 16'sd108, -16'sd76, 16'sd24, 16'sd75};
        weights1[37] = '{-16'sd20, 16'sd48, 16'sd169, 16'sd26, -16'sd97, 16'sd132, 16'sd108, -16'sd70, 16'sd84, -16'sd28, 16'sd20, -16'sd55, 16'sd28, -16'sd5, 16'sd175, -16'sd62, 16'sd52, 16'sd81, -16'sd5, 16'sd0, 16'sd59, -16'sd16, 16'sd13, 16'sd65, 16'sd123, -16'sd27, -16'sd69, 16'sd89, 16'sd132, -16'sd20, 16'sd11, 16'sd76};
        weights1[38] = '{-16'sd64, 16'sd6, 16'sd45, -16'sd69, -16'sd24, 16'sd164, -16'sd21, -16'sd58, 16'sd44, 16'sd44, -16'sd39, -16'sd38, 16'sd12, 16'sd40, 16'sd134, -16'sd83, -16'sd12, 16'sd105, 16'sd26, 16'sd72, 16'sd32, 16'sd8, -16'sd72, 16'sd4, -16'sd48, 16'sd79, -16'sd167, 16'sd88, 16'sd85, 16'sd10, 16'sd72, 16'sd115};
        weights1[39] = '{-16'sd176, -16'sd101, -16'sd262, -16'sd66, 16'sd78, 16'sd276, -16'sd101, 16'sd35, 16'sd76, -16'sd93, -16'sd169, 16'sd110, 16'sd80, 16'sd39, 16'sd150, -16'sd122, 16'sd195, 16'sd146, 16'sd153, 16'sd195, -16'sd121, -16'sd41, -16'sd54, -16'sd134, -16'sd60, 16'sd101, -16'sd246, 16'sd151, 16'sd53, 16'sd133, -16'sd27, -16'sd189};
        weights1[40] = '{-16'sd54, 16'sd120, 16'sd160, 16'sd28, -16'sd66, -16'sd132, -16'sd30, 16'sd173, -16'sd27, 16'sd237, 16'sd271, -16'sd8, 16'sd163, 16'sd100, -16'sd38, -16'sd194, 16'sd161, -16'sd236, 16'sd164, -16'sd263, 16'sd34, -16'sd112, 16'sd113, 16'sd162, 16'sd207, -16'sd63, -16'sd134, -16'sd141, 16'sd207, -16'sd226, -16'sd159, 16'sd76};
        weights1[41] = '{16'sd27, 16'sd41, -16'sd2, 16'sd71, 16'sd10, 16'sd27, 16'sd64, -16'sd89, -16'sd20, -16'sd159, -16'sd42, -16'sd21, -16'sd96, -16'sd10, 16'sd52, -16'sd93, -16'sd54, 16'sd35, 16'sd15, 16'sd61, 16'sd128, -16'sd34, 16'sd13, -16'sd76, -16'sd15, -16'sd82, -16'sd147, -16'sd58, 16'sd154, 16'sd13, 16'sd62, 16'sd4};
        weights1[42] = '{16'sd5, 16'sd14, -16'sd31, 16'sd38, 16'sd65, -16'sd16, 16'sd37, -16'sd66, 16'sd37, -16'sd123, -16'sd141, -16'sd39, -16'sd188, -16'sd20, 16'sd67, 16'sd87, -16'sd130, 16'sd165, -16'sd26, 16'sd106, 16'sd134, 16'sd25, 16'sd91, -16'sd16, -16'sd94, 16'sd38, 16'sd18, 16'sd19, 16'sd3, 16'sd60, 16'sd62, -16'sd79};
        weights1[43] = '{-16'sd9, -16'sd14, -16'sd17, 16'sd75, 16'sd69, 16'sd95, 16'sd86, -16'sd2, -16'sd63, -16'sd132, -16'sd22, -16'sd68, -16'sd53, 16'sd23, 16'sd24, 16'sd26, -16'sd79, -16'sd63, -16'sd88, 16'sd71, 16'sd57, 16'sd106, 16'sd20, -16'sd33, -16'sd111, -16'sd10, 16'sd86, 16'sd33, 16'sd74, 16'sd125, 16'sd56, -16'sd52};
        weights1[44] = '{-16'sd44, -16'sd21, -16'sd79, 16'sd63, 16'sd79, 16'sd37, 16'sd81, 16'sd46, 16'sd18, -16'sd144, -16'sd88, 16'sd1, -16'sd39, -16'sd95, 16'sd107, 16'sd65, 16'sd45, 16'sd38, -16'sd93, 16'sd84, -16'sd5, -16'sd11, -16'sd95, -16'sd185, -16'sd53, 16'sd14, 16'sd135, 16'sd63, 16'sd95, 16'sd76, -16'sd24, -16'sd17};
        weights1[45] = '{16'sd106, 16'sd85, -16'sd171, 16'sd85, -16'sd108, 16'sd17, 16'sd90, -16'sd10, 16'sd65, -16'sd64, 16'sd7, 16'sd16, -16'sd56, -16'sd125, 16'sd98, 16'sd142, 16'sd114, 16'sd70, -16'sd29, -16'sd74, -16'sd59, -16'sd57, 16'sd73, -16'sd121, 16'sd57, -16'sd84, -16'sd64, -16'sd25, -16'sd17, 16'sd68, 16'sd12, -16'sd72};
        weights1[46] = '{16'sd90, 16'sd44, 16'sd10, 16'sd91, -16'sd79, 16'sd11, 16'sd82, -16'sd55, -16'sd18, -16'sd100, -16'sd22, -16'sd43, -16'sd32, 16'sd38, 16'sd47, -16'sd37, -16'sd26, -16'sd36, 16'sd16, -16'sd68, 16'sd10, -16'sd11, 16'sd60, -16'sd7, -16'sd26, -16'sd31, 16'sd62, -16'sd17, 16'sd36, 16'sd16, 16'sd39, 16'sd72};
        weights1[47] = '{-16'sd4, 16'sd2, 16'sd31, 16'sd19, -16'sd87, 16'sd6, 16'sd42, -16'sd68, 16'sd42, -16'sd75, 16'sd71, 16'sd32, -16'sd82, -16'sd110, 16'sd22, -16'sd73, -16'sd70, 16'sd41, -16'sd91, -16'sd40, 16'sd116, 16'sd16, 16'sd41, -16'sd63, -16'sd10, -16'sd41, 16'sd64, 16'sd43, 16'sd15, -16'sd3, 16'sd33, 16'sd94};
        weights1[48] = '{-16'sd53, -16'sd81, 16'sd92, 16'sd26, -16'sd96, -16'sd91, 16'sd32, -16'sd73, 16'sd78, 16'sd21, 16'sd50, -16'sd37, -16'sd85, -16'sd116, 16'sd20, 16'sd51, -16'sd144, -16'sd102, -16'sd173, -16'sd59, 16'sd212, -16'sd25, -16'sd37, -16'sd61, -16'sd7, 16'sd103, 16'sd38, 16'sd124, 16'sd133, -16'sd63, 16'sd80, 16'sd23};
        weights1[49] = '{-16'sd117, -16'sd50, -16'sd178, -16'sd64, 16'sd59, 16'sd136, -16'sd140, -16'sd32, 16'sd25, 16'sd57, -16'sd52, 16'sd56, 16'sd149, 16'sd31, 16'sd0, -16'sd210, 16'sd297, 16'sd90, 16'sd165, 16'sd188, -16'sd271, -16'sd178, -16'sd33, -16'sd57, 16'sd154, 16'sd144, -16'sd184, 16'sd162, -16'sd36, -16'sd45, -16'sd115, 16'sd41};
        weights1[50] = '{16'sd11, 16'sd30, 16'sd45, -16'sd55, -16'sd24, -16'sd39, -16'sd52, 16'sd149, -16'sd117, 16'sd185, 16'sd168, 16'sd45, 16'sd229, 16'sd91, 16'sd45, -16'sd126, 16'sd194, -16'sd137, 16'sd102, -16'sd93, -16'sd143, -16'sd83, 16'sd30, 16'sd98, 16'sd161, -16'sd74, -16'sd164, -16'sd40, 16'sd57, -16'sd154, -16'sd201, 16'sd64};
        weights1[51] = '{-16'sd5, -16'sd44, 16'sd47, 16'sd38, 16'sd23, -16'sd69, -16'sd27, 16'sd147, -16'sd113, -16'sd60, -16'sd59, -16'sd52, -16'sd78, 16'sd20, 16'sd86, -16'sd157, 16'sd21, -16'sd10, -16'sd67, 16'sd40, -16'sd36, -16'sd50, 16'sd8, -16'sd123, 16'sd28, -16'sd81, -16'sd63, 16'sd97, -16'sd5, -16'sd42, 16'sd37, 16'sd129};
        weights1[52] = '{16'sd56, -16'sd19, 16'sd123, 16'sd9, 16'sd36, 16'sd11, -16'sd29, 16'sd49, -16'sd34, -16'sd24, 16'sd11, -16'sd15, -16'sd64, 16'sd42, 16'sd46, -16'sd51, -16'sd89, 16'sd71, -16'sd124, -16'sd7, 16'sd36, 16'sd65, -16'sd27, -16'sd101, -16'sd45, -16'sd37, 16'sd75, 16'sd89, 16'sd31, -16'sd33, 16'sd53, 16'sd2};
        weights1[53] = '{16'sd90, -16'sd88, 16'sd61, -16'sd35, 16'sd60, 16'sd94, 16'sd29, 16'sd138, 16'sd2, 16'sd38, -16'sd50, 16'sd7, 16'sd23, 16'sd21, 16'sd65, -16'sd85, -16'sd87, 16'sd16, -16'sd80, 16'sd61, 16'sd98, 16'sd5, -16'sd15, -16'sd82, 16'sd6, -16'sd8, 16'sd113, 16'sd100, -16'sd24, 16'sd33, 16'sd59, 16'sd26};
        weights1[54] = '{16'sd103, -16'sd66, -16'sd17, 16'sd26, -16'sd99, 16'sd30, 16'sd123, 16'sd13, 16'sd96, -16'sd32, 16'sd131, 16'sd9, 16'sd114, 16'sd47, -16'sd30, 16'sd48, 16'sd101, 16'sd8, 16'sd3, 16'sd86, -16'sd44, 16'sd70, -16'sd103, -16'sd126, 16'sd108, 16'sd52, 16'sd144, 16'sd10, -16'sd40, 16'sd97, -16'sd11, 16'sd7};
        weights1[55] = '{16'sd121, -16'sd37, -16'sd120, -16'sd38, -16'sd81, 16'sd89, 16'sd131, 16'sd3, 16'sd31, -16'sd83, 16'sd86, 16'sd49, 16'sd35, -16'sd1, 16'sd55, 16'sd60, 16'sd37, 16'sd5, -16'sd23, -16'sd167, -16'sd43, 16'sd4, 16'sd65, -16'sd66, 16'sd41, -16'sd24, 16'sd7, -16'sd108, -16'sd107, 16'sd45, 16'sd14, -16'sd131};
        weights1[56] = '{16'sd23, 16'sd58, -16'sd37, 16'sd90, -16'sd27, 16'sd67, 16'sd65, 16'sd52, -16'sd65, 16'sd45, 16'sd0, 16'sd4, 16'sd44, 16'sd70, 16'sd82, 16'sd15, -16'sd16, -16'sd127, -16'sd55, -16'sd103, 16'sd36, 16'sd102, 16'sd40, -16'sd107, -16'sd12, -16'sd15, 16'sd74, 16'sd63, 16'sd38, 16'sd81, 16'sd11, 16'sd91};
        weights1[57] = '{16'sd11, 16'sd108, -16'sd24, 16'sd55, 16'sd101, -16'sd135, 16'sd66, 16'sd64, -16'sd112, 16'sd42, -16'sd69, -16'sd41, -16'sd9, 16'sd32, 16'sd7, 16'sd28, -16'sd30, -16'sd1, 16'sd25, -16'sd28, 16'sd73, 16'sd34, 16'sd21, -16'sd56, 16'sd61, -16'sd53, 16'sd42, 16'sd89, 16'sd77, 16'sd0, -16'sd15, -16'sd55};
        weights1[58] = '{-16'sd49, 16'sd31, 16'sd19, 16'sd0, 16'sd99, -16'sd156, 16'sd23, 16'sd87, -16'sd44, 16'sd126, -16'sd114, 16'sd29, 16'sd31, 16'sd93, 16'sd34, 16'sd20, -16'sd59, 16'sd31, -16'sd60, 16'sd9, 16'sd77, -16'sd17, 16'sd36, 16'sd2, 16'sd17, 16'sd5, 16'sd60, 16'sd58, 16'sd171, -16'sd3, -16'sd124, -16'sd44};
        weights1[59] = '{16'sd167, -16'sd72, -16'sd115, 16'sd22, -16'sd207, -16'sd67, -16'sd61, 16'sd13, 16'sd56, 16'sd235, 16'sd122, 16'sd121, 16'sd201, -16'sd27, -16'sd169, -16'sd129, 16'sd89, -16'sd43, -16'sd62, -16'sd101, -16'sd174, -16'sd149, 16'sd4, 16'sd21, 16'sd130, 16'sd72, 16'sd49, 16'sd25, -16'sd107, -16'sd120, -16'sd207, 16'sd67};
        weights1[60] = '{-16'sd17, -16'sd17, -16'sd134, -16'sd67, 16'sd173, 16'sd140, 16'sd24, 16'sd196, -16'sd193, -16'sd99, -16'sd198, 16'sd25, 16'sd123, 16'sd172, 16'sd220, -16'sd128, 16'sd222, 16'sd116, 16'sd149, 16'sd255, -16'sd255, -16'sd130, -16'sd28, -16'sd68, 16'sd45, 16'sd25, -16'sd131, 16'sd119, -16'sd66, 16'sd141, -16'sd118, -16'sd50};
        weights1[61] = '{16'sd57, -16'sd3, 16'sd40, 16'sd4, 16'sd7, -16'sd85, 16'sd8, 16'sd137, -16'sd138, -16'sd5, 16'sd0, 16'sd44, 16'sd132, 16'sd55, 16'sd72, -16'sd174, 16'sd128, -16'sd77, 16'sd68, 16'sd128, -16'sd214, -16'sd41, -16'sd24, -16'sd14, 16'sd41, 16'sd56, -16'sd87, 16'sd122, -16'sd50, -16'sd54, -16'sd104, 16'sd105};
        weights1[62] = '{16'sd53, 16'sd23, 16'sd34, -16'sd55, -16'sd60, 16'sd22, 16'sd32, 16'sd78, -16'sd5, 16'sd37, -16'sd2, 16'sd4, -16'sd10, 16'sd50, 16'sd38, -16'sd37, -16'sd55, 16'sd13, -16'sd140, 16'sd29, -16'sd76, -16'sd15, -16'sd130, -16'sd48, 16'sd54, 16'sd43, -16'sd19, 16'sd130, -16'sd40, -16'sd3, -16'sd23, 16'sd97};
        weights1[63] = '{-16'sd18, 16'sd53, 16'sd59, -16'sd17, -16'sd54, -16'sd62, 16'sd15, -16'sd66, 16'sd103, 16'sd88, 16'sd25, 16'sd100, -16'sd80, -16'sd95, 16'sd19, -16'sd39, -16'sd94, 16'sd21, -16'sd122, -16'sd26, 16'sd69, 16'sd86, -16'sd93, 16'sd8, 16'sd27, 16'sd75, 16'sd110, 16'sd26, 16'sd38, -16'sd56, 16'sd26, 16'sd2};
        weights1[64] = '{16'sd53, 16'sd16, -16'sd32, -16'sd57, -16'sd119, 16'sd32, 16'sd41, 16'sd37, 16'sd117, 16'sd58, 16'sd125, 16'sd94, -16'sd23, 16'sd48, -16'sd83, 16'sd87, 16'sd85, 16'sd180, 16'sd4, -16'sd119, 16'sd133, 16'sd64, 16'sd8, -16'sd29, 16'sd55, 16'sd130, 16'sd2, 16'sd7, -16'sd19, -16'sd63, -16'sd26, -16'sd54};
        weights1[65] = '{16'sd92, 16'sd36, -16'sd34, -16'sd5, -16'sd64, 16'sd141, 16'sd4, 16'sd113, -16'sd29, 16'sd68, 16'sd43, 16'sd33, -16'sd45, 16'sd131, -16'sd24, 16'sd101, 16'sd125, -16'sd88, -16'sd18, -16'sd74, 16'sd9, 16'sd98, 16'sd39, -16'sd88, 16'sd25, 16'sd3, 16'sd13, 16'sd86, -16'sd75, -16'sd25, 16'sd48, -16'sd87};
        weights1[66] = '{16'sd23, 16'sd29, 16'sd90, 16'sd38, 16'sd70, -16'sd34, 16'sd101, 16'sd109, -16'sd49, 16'sd35, -16'sd34, 16'sd91, 16'sd34, 16'sd84, 16'sd9, -16'sd34, -16'sd25, -16'sd118, 16'sd35, 16'sd9, 16'sd32, -16'sd7, -16'sd11, -16'sd80, 16'sd83, 16'sd20, 16'sd14, 16'sd94, 16'sd61, 16'sd97, 16'sd28, 16'sd28};
        weights1[67] = '{16'sd66, -16'sd7, 16'sd39, 16'sd29, 16'sd83, -16'sd86, 16'sd78, 16'sd49, -16'sd35, 16'sd29, 16'sd7, 16'sd12, 16'sd26, 16'sd18, 16'sd16, -16'sd40, 16'sd77, 16'sd21, 16'sd104, 16'sd14, -16'sd14, 16'sd3, -16'sd33, 16'sd9, 16'sd25, 16'sd42, 16'sd45, 16'sd46, -16'sd3, 16'sd5, -16'sd4, -16'sd69};
        weights1[68] = '{16'sd78, 16'sd3, -16'sd14, -16'sd11, 16'sd65, -16'sd161, -16'sd2, 16'sd56, 16'sd59, 16'sd69, 16'sd76, 16'sd84, 16'sd81, 16'sd8, -16'sd40, -16'sd80, 16'sd23, 16'sd35, 16'sd36, 16'sd103, -16'sd68, -16'sd75, 16'sd8, 16'sd0, 16'sd27, 16'sd19, 16'sd61, 16'sd89, 16'sd130, -16'sd29, -16'sd52, -16'sd11};
        weights1[69] = '{16'sd118, -16'sd96, 16'sd109, -16'sd21, -16'sd109, -16'sd129, -16'sd107, 16'sd166, 16'sd107, 16'sd238, 16'sd139, 16'sd125, 16'sd149, 16'sd76, -16'sd141, -16'sd123, -16'sd47, 16'sd81, -16'sd83, -16'sd226, -16'sd89, -16'sd127, 16'sd56, 16'sd58, 16'sd157, 16'sd56, 16'sd198, -16'sd9, -16'sd217, -16'sd235, -16'sd138, 16'sd98};
        weights1[70] = '{-16'sd42, -16'sd76, -16'sd138, -16'sd35, 16'sd178, 16'sd62, 16'sd31, 16'sd170, -16'sd200, -16'sd15, -16'sd115, -16'sd5, 16'sd88, 16'sd262, 16'sd156, -16'sd81, 16'sd198, 16'sd113, 16'sd180, 16'sd197, -16'sd267, -16'sd14, -16'sd85, -16'sd111, -16'sd11, 16'sd72, -16'sd120, 16'sd142, 16'sd15, 16'sd194, -16'sd46, 16'sd35};
        weights1[71] = '{16'sd35, -16'sd37, 16'sd33, -16'sd11, -16'sd31, 16'sd18, -16'sd3, 16'sd11, -16'sd19, 16'sd70, 16'sd59, 16'sd38, 16'sd81, 16'sd86, 16'sd41, -16'sd144, 16'sd106, -16'sd116, 16'sd87, 16'sd80, -16'sd132, -16'sd94, -16'sd9, -16'sd22, 16'sd83, -16'sd11, 16'sd21, 16'sd77, -16'sd88, -16'sd19, -16'sd47, 16'sd55};
        weights1[72] = '{-16'sd3, -16'sd12, 16'sd70, -16'sd24, -16'sd44, 16'sd2, -16'sd3, -16'sd79, 16'sd68, 16'sd28, 16'sd34, 16'sd77, 16'sd51, -16'sd14, 16'sd50, -16'sd34, 16'sd32, -16'sd101, 16'sd127, 16'sd82, -16'sd123, -16'sd75, -16'sd42, -16'sd12, 16'sd88, 16'sd91, -16'sd69, 16'sd77, -16'sd15, -16'sd128, 16'sd41, 16'sd35};
        weights1[73] = '{16'sd0, -16'sd53, 16'sd104, -16'sd95, 16'sd20, -16'sd111, 16'sd35, -16'sd9, 16'sd81, 16'sd76, 16'sd15, 16'sd49, 16'sd22, 16'sd17, 16'sd53, -16'sd2, 16'sd48, 16'sd72, -16'sd13, 16'sd76, 16'sd52, -16'sd61, -16'sd55, 16'sd25, 16'sd57, 16'sd51, -16'sd68, 16'sd96, 16'sd56, -16'sd110, -16'sd86, 16'sd34};
        weights1[74] = '{-16'sd18, -16'sd25, 16'sd15, -16'sd86, 16'sd75, -16'sd102, 16'sd38, 16'sd55, -16'sd6, 16'sd87, 16'sd19, 16'sd84, -16'sd72, 16'sd31, 16'sd17, 16'sd69, -16'sd29, 16'sd93, 16'sd7, 16'sd56, 16'sd70, 16'sd3, -16'sd33, 16'sd82, 16'sd43, 16'sd88, 16'sd4, 16'sd28, 16'sd174, -16'sd54, 16'sd37, -16'sd42};
        weights1[75] = '{16'sd84, -16'sd63, -16'sd24, -16'sd112, 16'sd68, -16'sd79, 16'sd87, 16'sd62, -16'sd4, -16'sd12, -16'sd30, 16'sd31, -16'sd66, -16'sd12, -16'sd10, 16'sd92, 16'sd63, -16'sd232, 16'sd100, 16'sd107, 16'sd27, -16'sd5, 16'sd54, 16'sd70, 16'sd48, 16'sd56, -16'sd2, 16'sd40, 16'sd53, -16'sd23, -16'sd12, 16'sd14};
        weights1[76] = '{16'sd127, -16'sd115, 16'sd63, 16'sd19, 16'sd32, -16'sd55, -16'sd23, 16'sd9, 16'sd25, -16'sd65, 16'sd13, 16'sd99, 16'sd20, 16'sd9, 16'sd16, 16'sd49, 16'sd24, -16'sd59, 16'sd93, 16'sd34, 16'sd1, 16'sd32, -16'sd43, 16'sd54, 16'sd39, 16'sd46, -16'sd22, -16'sd20, 16'sd45, 16'sd75, -16'sd73, 16'sd51};
        weights1[77] = '{16'sd105, -16'sd66, -16'sd2, 16'sd15, 16'sd20, -16'sd130, 16'sd7, -16'sd73, 16'sd105, 16'sd49, 16'sd30, 16'sd17, -16'sd2, -16'sd60, -16'sd41, -16'sd80, 16'sd55, 16'sd14, 16'sd8, 16'sd40, -16'sd95, -16'sd42, -16'sd46, 16'sd25, -16'sd3, 16'sd68, -16'sd45, 16'sd47, -16'sd45, 16'sd37, -16'sd45, 16'sd2};
        weights1[78] = '{16'sd92, -16'sd61, -16'sd57, -16'sd36, 16'sd19, -16'sd121, -16'sd132, -16'sd100, 16'sd156, 16'sd60, 16'sd29, 16'sd47, 16'sd38, 16'sd51, -16'sd77, -16'sd140, -16'sd22, 16'sd100, -16'sd12, 16'sd52, -16'sd68, 16'sd9, -16'sd54, -16'sd26, 16'sd21, 16'sd69, -16'sd58, 16'sd135, -16'sd22, -16'sd64, 16'sd0, -16'sd9};
        weights1[79] = '{16'sd27, -16'sd26, 16'sd1, -16'sd78, -16'sd98, -16'sd96, -16'sd190, 16'sd34, 16'sd89, 16'sd127, 16'sd148, 16'sd55, 16'sd125, 16'sd107, -16'sd136, -16'sd93, -16'sd79, 16'sd72, -16'sd175, -16'sd114, -16'sd177, -16'sd98, -16'sd3, 16'sd114, 16'sd120, 16'sd95, 16'sd4, 16'sd21, -16'sd136, -16'sd129, -16'sd29, 16'sd33};
        weights1[80] = '{-16'sd15, -16'sd12, -16'sd174, -16'sd90, 16'sd141, 16'sd133, 16'sd39, 16'sd137, -16'sd125, -16'sd79, -16'sd239, -16'sd22, 16'sd59, 16'sd160, 16'sd192, -16'sd73, 16'sd198, 16'sd158, 16'sd144, 16'sd248, -16'sd298, -16'sd61, -16'sd5, -16'sd46, 16'sd22, 16'sd25, -16'sd172, 16'sd171, -16'sd54, 16'sd256, -16'sd57, -16'sd4};
        weights1[81] = '{16'sd23, 16'sd43, -16'sd6, 16'sd10, 16'sd36, 16'sd22, -16'sd48, 16'sd88, -16'sd56, 16'sd46, -16'sd2, 16'sd62, 16'sd120, 16'sd80, 16'sd94, -16'sd26, 16'sd154, 16'sd52, 16'sd71, 16'sd67, -16'sd108, -16'sd74, 16'sd54, 16'sd64, 16'sd73, -16'sd22, -16'sd49, -16'sd58, -16'sd10, 16'sd82, -16'sd87, -16'sd34};
        weights1[82] = '{16'sd7, 16'sd44, 16'sd113, 16'sd64, 16'sd4, 16'sd31, 16'sd22, 16'sd0, 16'sd14, -16'sd51, 16'sd43, 16'sd18, 16'sd74, -16'sd13, 16'sd38, -16'sd9, 16'sd40, 16'sd45, 16'sd35, -16'sd10, 16'sd30, -16'sd51, -16'sd25, 16'sd75, 16'sd36, -16'sd42, -16'sd2, -16'sd58, -16'sd36, -16'sd12, -16'sd11, 16'sd56};
        weights1[83] = '{16'sd10, -16'sd1, 16'sd98, 16'sd18, 16'sd66, 16'sd49, 16'sd90, 16'sd13, 16'sd24, -16'sd48, 16'sd46, 16'sd16, 16'sd77, 16'sd27, 16'sd18, -16'sd20, -16'sd8, 16'sd34, 16'sd65, 16'sd32, -16'sd3, 16'sd54, -16'sd3, 16'sd44, 16'sd3, -16'sd1, -16'sd59, 16'sd36, 16'sd58, -16'sd7, 16'sd48, 16'sd38};
        weights1[84] = '{16'sd38, 16'sd45, 16'sd27, 16'sd45, 16'sd39, -16'sd1, 16'sd112, -16'sd22, 16'sd118, 16'sd33, -16'sd25, 16'sd77, 16'sd100, 16'sd25, 16'sd100, 16'sd7, 16'sd80, 16'sd37, 16'sd72, 16'sd46, 16'sd107, 16'sd79, 16'sd25, 16'sd59, -16'sd20, 16'sd63, -16'sd40, 16'sd26, 16'sd87, 16'sd19, 16'sd19, 16'sd87};
        weights1[85] = '{16'sd41, 16'sd41, -16'sd17, 16'sd3, 16'sd69, 16'sd25, 16'sd17, -16'sd99, 16'sd39, -16'sd24, 16'sd33, 16'sd66, 16'sd22, 16'sd83, 16'sd114, 16'sd121, 16'sd41, -16'sd131, 16'sd37, 16'sd65, 16'sd65, 16'sd80, -16'sd2, 16'sd61, -16'sd17, 16'sd71, -16'sd49, -16'sd23, 16'sd108, 16'sd23, -16'sd20, 16'sd40};
        weights1[86] = '{16'sd96, -16'sd112, 16'sd37, 16'sd3, 16'sd19, -16'sd40, -16'sd29, -16'sd44, 16'sd96, -16'sd65, -16'sd28, 16'sd7, 16'sd56, -16'sd28, -16'sd14, 16'sd24, 16'sd90, -16'sd47, 16'sd68, 16'sd19, 16'sd4, 16'sd124, 16'sd0, 16'sd92, 16'sd62, 16'sd12, -16'sd34, -16'sd31, 16'sd12, 16'sd81, 16'sd57, -16'sd28};
        weights1[87] = '{16'sd125, -16'sd132, -16'sd8, 16'sd2, 16'sd35, -16'sd50, 16'sd44, -16'sd88, 16'sd94, 16'sd18, 16'sd66, 16'sd52, 16'sd41, 16'sd24, -16'sd61, -16'sd62, -16'sd49, 16'sd83, -16'sd5, 16'sd15, -16'sd88, 16'sd78, -16'sd107, -16'sd4, 16'sd77, 16'sd33, 16'sd40, 16'sd17, -16'sd38, 16'sd71, 16'sd84, 16'sd15};
        weights1[88] = '{16'sd91, -16'sd91, 16'sd24, 16'sd30, -16'sd21, 16'sd2, 16'sd21, -16'sd76, 16'sd84, -16'sd11, 16'sd21, 16'sd61, 16'sd71, 16'sd45, -16'sd97, -16'sd159, -16'sd133, 16'sd153, 16'sd17, 16'sd41, -16'sd107, 16'sd129, -16'sd40, 16'sd3, 16'sd28, 16'sd55, -16'sd86, 16'sd93, -16'sd59, -16'sd3, 16'sd109, 16'sd35};
        weights1[89] = '{16'sd41, -16'sd125, -16'sd3, -16'sd65, -16'sd70, -16'sd155, -16'sd161, 16'sd134, -16'sd29, 16'sd173, 16'sd99, 16'sd106, 16'sd184, 16'sd93, -16'sd163, -16'sd102, -16'sd23, 16'sd102, -16'sd189, -16'sd78, -16'sd182, -16'sd48, -16'sd10, 16'sd95, 16'sd55, 16'sd90, -16'sd78, 16'sd106, -16'sd143, -16'sd115, -16'sd57, 16'sd51};
        weights1[90] = '{16'sd49, 16'sd124, 16'sd6, 16'sd125, 16'sd155, 16'sd138, 16'sd178, 16'sd98, -16'sd178, -16'sd57, -16'sd176, -16'sd111, 16'sd151, 16'sd70, 16'sd201, -16'sd19, 16'sd156, 16'sd80, 16'sd149, 16'sd12, -16'sd22, -16'sd84, 16'sd51, 16'sd170, 16'sd3, -16'sd192, -16'sd135, -16'sd167, 16'sd111, 16'sd173, -16'sd141, 16'sd87};
        weights1[91] = '{16'sd2, 16'sd116, 16'sd88, 16'sd115, 16'sd29, 16'sd69, 16'sd172, 16'sd17, -16'sd98, 16'sd7, -16'sd202, -16'sd60, 16'sd18, 16'sd11, 16'sd101, -16'sd46, 16'sd82, 16'sd89, 16'sd46, -16'sd3, 16'sd91, 16'sd44, 16'sd151, 16'sd144, -16'sd41, -16'sd139, -16'sd158, -16'sd119, -16'sd2, 16'sd172, 16'sd9, 16'sd166};
        weights1[92] = '{16'sd4, 16'sd92, 16'sd66, 16'sd180, 16'sd5, 16'sd53, 16'sd148, -16'sd60, -16'sd39, -16'sd63, -16'sd110, 16'sd13, 16'sd191, 16'sd5, 16'sd111, -16'sd46, 16'sd80, 16'sd9, 16'sd102, -16'sd45, -16'sd7, -16'sd98, 16'sd49, 16'sd83, -16'sd21, -16'sd102, -16'sd203, -16'sd121, 16'sd61, 16'sd102, 16'sd85, 16'sd105};
        weights1[93] = '{16'sd83, 16'sd41, -16'sd153, 16'sd87, 16'sd45, 16'sd54, 16'sd153, -16'sd111, -16'sd75, -16'sd10, -16'sd58, -16'sd38, 16'sd184, -16'sd8, 16'sd61, -16'sd98, 16'sd52, -16'sd19, 16'sd142, 16'sd82, -16'sd14, -16'sd60, 16'sd72, 16'sd89, 16'sd52, -16'sd142, -16'sd172, -16'sd71, -16'sd35, 16'sd125, 16'sd33, 16'sd159};
        weights1[94] = '{16'sd26, 16'sd100, -16'sd144, 16'sd70, 16'sd70, 16'sd59, 16'sd126, -16'sd102, -16'sd65, 16'sd40, -16'sd56, -16'sd12, 16'sd176, -16'sd9, -16'sd7, -16'sd107, 16'sd33, -16'sd31, 16'sd198, 16'sd110, -16'sd14, -16'sd129, 16'sd89, 16'sd57, 16'sd35, -16'sd99, -16'sd117, -16'sd22, -16'sd95, 16'sd130, 16'sd55, 16'sd130};
        weights1[95] = '{-16'sd19, 16'sd141, -16'sd170, 16'sd50, 16'sd40, 16'sd88, 16'sd70, -16'sd110, -16'sd23, 16'sd63, -16'sd17, -16'sd51, 16'sd165, 16'sd38, 16'sd36, -16'sd119, 16'sd25, -16'sd102, 16'sd208, 16'sd75, 16'sd42, -16'sd62, 16'sd108, 16'sd41, -16'sd86, 16'sd9, -16'sd149, -16'sd61, -16'sd105, 16'sd116, 16'sd86, 16'sd143};
        weights1[96] = '{-16'sd87, 16'sd174, -16'sd104, 16'sd112, 16'sd37, 16'sd121, 16'sd67, -16'sd173, -16'sd105, 16'sd28, -16'sd74, -16'sd32, 16'sd117, -16'sd82, 16'sd41, -16'sd181, -16'sd41, -16'sd95, 16'sd230, 16'sd83, 16'sd64, -16'sd45, 16'sd70, 16'sd59, -16'sd55, 16'sd30, -16'sd149, -16'sd68, -16'sd64, -16'sd9, 16'sd106, 16'sd110};
        weights1[97] = '{-16'sd20, 16'sd169, -16'sd120, 16'sd147, -16'sd16, 16'sd109, 16'sd57, -16'sd118, -16'sd22, -16'sd109, -16'sd95, -16'sd76, 16'sd77, -16'sd84, 16'sd24, -16'sd163, -16'sd145, 16'sd0, 16'sd73, 16'sd42, 16'sd134, -16'sd14, 16'sd90, -16'sd40, -16'sd105, -16'sd85, -16'sd165, -16'sd96, -16'sd16, 16'sd102, 16'sd76, 16'sd147};
        weights1[98] = '{-16'sd19, 16'sd55, -16'sd65, 16'sd67, 16'sd113, 16'sd98, 16'sd4, -16'sd50, -16'sd13, -16'sd129, -16'sd172, 16'sd25, -16'sd42, 16'sd10, 16'sd111, -16'sd9, -16'sd6, 16'sd47, 16'sd0, 16'sd45, -16'sd11, 16'sd32, -16'sd31, -16'sd26, -16'sd162, 16'sd55, -16'sd84, -16'sd47, -16'sd26, 16'sd144, 16'sd17, -16'sd7};
        weights1[99] = '{16'sd79, -16'sd36, -16'sd52, -16'sd65, -16'sd3, -16'sd18, -16'sd72, -16'sd7, 16'sd46, 16'sd41, 16'sd55, 16'sd89, 16'sd96, -16'sd14, -16'sd134, -16'sd88, -16'sd73, -16'sd25, -16'sd8, 16'sd21, -16'sd83, 16'sd1, -16'sd3, 16'sd74, 16'sd31, 16'sd32, -16'sd6, 16'sd21, -16'sd85, -16'sd58, -16'sd27, 16'sd31};

    end

    logic signed [15:0] weights2 [32][16];
    initial begin  
        weights2[0] = '{16'sd7, 16'sd125, 16'sd49, 16'sd136, 16'sd79, -16'sd133, -16'sd30, -16'sd60, 16'sd62, 16'sd122, 16'sd125, -16'sd80, 16'sd80, 16'sd98, 16'sd113, 16'sd5};
        weights2[1] = '{16'sd171, 16'sd122, 16'sd25, -16'sd160, -16'sd129, 16'sd155, -16'sd86, -16'sd28, -16'sd103, 16'sd8, -16'sd101, -16'sd27, 16'sd58, 16'sd13, -16'sd97, -16'sd46};
        weights2[2] = '{16'sd78, -16'sd156, -16'sd78, 16'sd120, 16'sd16, 16'sd18, -16'sd164, 16'sd95, 16'sd2, -16'sd154, 16'sd8, 16'sd24, -16'sd169, 16'sd53, -16'sd180, 16'sd132};
        weights2[3] = '{16'sd143, 16'sd103, 16'sd122, 16'sd83, 16'sd190, -16'sd273, 16'sd53, -16'sd151, 16'sd91, 16'sd149, -16'sd156, 16'sd30, 16'sd82, 16'sd161, -16'sd249, -16'sd95};
        weights2[4] = '{16'sd162, 16'sd167, -16'sd103, -16'sd73, 16'sd17, 16'sd6, -16'sd116, -16'sd138, -16'sd151, -16'sd50, -16'sd75, 16'sd54, 16'sd42, 16'sd135, 16'sd6, -16'sd49};
        weights2[5] = '{16'sd111, 16'sd85, -16'sd39, 16'sd98, -16'sd164, 16'sd200, -16'sd78, -16'sd26, -16'sd128, 16'sd88, 16'sd174, 16'sd131, 16'sd13, 16'sd4, 16'sd11, -16'sd99};
        weights2[6] = '{-16'sd2, 16'sd139, -16'sd43, 16'sd122, 16'sd80, 16'sd76, 16'sd49, 16'sd48, 16'sd5, 16'sd82, 16'sd1, -16'sd78, 16'sd26, 16'sd106, 16'sd100, 16'sd152};
        weights2[7] = '{16'sd52, -16'sd146, 16'sd218, 16'sd150, 16'sd82, -16'sd59, -16'sd25, 16'sd40, -16'sd14, -16'sd90, 16'sd35, -16'sd98, -16'sd71, 16'sd9, -16'sd202, 16'sd165};
        weights2[8] = '{-16'sd79, 16'sd159, 16'sd15, -16'sd80, -16'sd44, -16'sd71, 16'sd179, 16'sd40, 16'sd153, 16'sd49, 16'sd122, 16'sd60, -16'sd90, -16'sd182, 16'sd157, -16'sd80};
        weights2[9] = '{16'sd93, -16'sd223, 16'sd166, 16'sd15, 16'sd105, 16'sd138, 16'sd18, -16'sd157, 16'sd32, 16'sd2, -16'sd130, 16'sd58, 16'sd121, 16'sd39, 16'sd62, 16'sd74};
        weights2[10] = '{-16'sd42, 16'sd154, 16'sd211, -16'sd44, 16'sd124, -16'sd110, 16'sd145, 16'sd16, 16'sd118, 16'sd14, -16'sd84, 16'sd57, 16'sd168, -16'sd75, 16'sd40, -16'sd56};
        weights2[11] = '{-16'sd105, 16'sd103, 16'sd33, 16'sd12, 16'sd77, -16'sd116, 16'sd27, 16'sd111, 16'sd108, -16'sd34, 16'sd117, -16'sd1, 16'sd35, -16'sd111, 16'sd82, 16'sd90};
        weights2[12] = '{-16'sd29, 16'sd161, 16'sd172, 16'sd53, -16'sd60, 16'sd132, -16'sd71, -16'sd110, 16'sd83, -16'sd115, -16'sd35, 16'sd85, 16'sd40, -16'sd50, 16'sd85, 16'sd129};
        weights2[13] = '{16'sd141, -16'sd129, 16'sd186, 16'sd142, 16'sd55, 16'sd153, -16'sd49, -16'sd31, -16'sd5, 16'sd106, 16'sd75, 16'sd44, 16'sd21, 16'sd50, 16'sd92, 16'sd90};
        weights2[14] = '{16'sd55, 16'sd73, -16'sd48, -16'sd7, -16'sd133, 16'sd104, -16'sd18, -16'sd44, 16'sd45, 16'sd112, 16'sd131, 16'sd50, -16'sd101, 16'sd44, -16'sd49, 16'sd40};
        weights2[15] = '{-16'sd111, 16'sd22, -16'sd33, 16'sd35, -16'sd56, -16'sd58, 16'sd204, 16'sd171, -16'sd31, 16'sd81, 16'sd148, -16'sd104, 16'sd118, 16'sd104, -16'sd66, -16'sd47};
        weights2[16] = '{16'sd68, 16'sd146, 16'sd154, 16'sd32, -16'sd137, 16'sd37, 16'sd91, 16'sd7, 16'sd6, -16'sd137, 16'sd165, 16'sd7, -16'sd79, -16'sd9, -16'sd82, 16'sd17};
        weights2[17] = '{16'sd193, -16'sd225, 16'sd41, -16'sd39, -16'sd147, 16'sd12, -16'sd12, 16'sd319, -16'sd81, -16'sd110, 16'sd231, 16'sd235, 16'sd43, 16'sd125, -16'sd159, -16'sd169};
        weights2[18] = '{-16'sd7, 16'sd103, 16'sd91, -16'sd116, -16'sd150, 16'sd92, -16'sd75, 16'sd83, 16'sd78, -16'sd169, 16'sd84, 16'sd20, 16'sd48, -16'sd147, -16'sd51, 16'sd130};
        weights2[19] = '{16'sd45, -16'sd1, -16'sd191, 16'sd6, -16'sd23, 16'sd73, -16'sd151, 16'sd103, 16'sd103, -16'sd166, 16'sd36, 16'sd186, -16'sd174, -16'sd141, 16'sd58, 16'sd51};
        weights2[20] = '{16'sd109, -16'sd11, -16'sd152, -16'sd24, 16'sd160, 16'sd155, 16'sd117, 16'sd35, 16'sd90, 16'sd215, -16'sd188, -16'sd43, 16'sd93, 16'sd0, 16'sd5, 16'sd37};
        weights2[21] = '{16'sd134, -16'sd80, -16'sd25, 16'sd64, 16'sd105, 16'sd44, 16'sd113, -16'sd29, -16'sd25, 16'sd134, 16'sd137, 16'sd104, -16'sd4, 16'sd111, 16'sd121, 16'sd0};
        weights2[22] = '{16'sd150, 16'sd125, 16'sd47, -16'sd112, -16'sd27, 16'sd66, 16'sd18, 16'sd105, -16'sd85, -16'sd137, -16'sd130, -16'sd28, 16'sd214, 16'sd153, -16'sd115, -16'sd95};
        weights2[23] = '{16'sd130, -16'sd199, 16'sd256, 16'sd56, -16'sd124, -16'sd34, 16'sd106, -16'sd232, 16'sd91, -16'sd75, -16'sd19, 16'sd59, 16'sd54, -16'sd179, -16'sd188, 16'sd164};
        weights2[24] = '{-16'sd135, 16'sd87, 16'sd130, -16'sd19, 16'sd95, -16'sd49, -16'sd54, -16'sd87, 16'sd81, -16'sd86, 16'sd3, -16'sd81, 16'sd24, -16'sd83, -16'sd31, 16'sd43};
        weights2[25] = '{-16'sd150, -16'sd95, 16'sd41, 16'sd23, -16'sd13, 16'sd45, 16'sd36, 16'sd110, 16'sd132, 16'sd38, 16'sd0, 16'sd102, -16'sd79, -16'sd206, 16'sd92, 16'sd36};
        weights2[26] = '{16'sd26, -16'sd191, -16'sd4, 16'sd129, 16'sd214, -16'sd244, 16'sd85, 16'sd42, 16'sd91, 16'sd50, -16'sd135, 16'sd99, -16'sd49, 16'sd30, 16'sd23, -16'sd6};
        weights2[27] = '{-16'sd56, -16'sd97, -16'sd6, 16'sd1, 16'sd72, 16'sd117, -16'sd134, 16'sd59, 16'sd138, 16'sd72, 16'sd73, 16'sd131, -16'sd89, 16'sd50, 16'sd44, 16'sd94};
        weights2[28] = '{16'sd59, -16'sd39, -16'sd138, 16'sd26, -16'sd7, 16'sd80, 16'sd75, -16'sd101, 16'sd84, 16'sd33, -16'sd16, -16'sd60, 16'sd4, -16'sd106, -16'sd67, 16'sd154};
        weights2[29] = '{16'sd15, 16'sd15, -16'sd73, 16'sd125, -16'sd133, 16'sd91, 16'sd6, 16'sd129, -16'sd162, 16'sd35, 16'sd162, -16'sd66, -16'sd62, 16'sd136, 16'sd151, 16'sd56};
        weights2[30] = '{16'sd121, 16'sd65, -16'sd106, -16'sd41, 16'sd104, 16'sd98, -16'sd65, 16'sd119, 16'sd37, 16'sd66, -16'sd38, 16'sd129, 16'sd86, 16'sd91, 16'sd114, -16'sd132};
        weights2[31] = '{16'sd109, 16'sd149, 16'sd15, -16'sd42, 16'sd151, 16'sd92, -16'sd165, -16'sd141, 16'sd151, -16'sd36, -16'sd162, 16'sd45, -16'sd28, 16'sd35, 16'sd67, 16'sd54};
    end

    logic signed [15:0] weights3 [16][10];
    initial begin
        weights3[0] = '{16'sd140, -16'sd154, -16'sd99, -16'sd50, 16'sd49, -16'sd17, -16'sd205, 16'sd202, -16'sd141, 16'sd69};
        weights3[1] = '{-16'sd116, 16'sd75, -16'sd62, 16'sd184, -16'sd161, -16'sd163, -16'sd230, -16'sd49, 16'sd123, 16'sd110};
        weights3[2] = '{-16'sd188, 16'sd94, 16'sd205, 16'sd7, -16'sd78, -16'sd48, -16'sd177, 16'sd153, -16'sd229, -16'sd288};
        weights3[3] = '{-16'sd29, -16'sd127, -16'sd36, 16'sd76, 16'sd197, 16'sd9, 16'sd42, -16'sd171, -16'sd208, -16'sd180};
        weights3[4] = '{16'sd58, -16'sd210, 16'sd70, -16'sd65, 16'sd47, -16'sd185, 16'sd112, -16'sd100, -16'sd132, 16'sd92};
        weights3[5] = '{-16'sd11, -16'sd223, -16'sd119, 16'sd53, -16'sd66, 16'sd197, -16'sd86, 16'sd107, 16'sd59, -16'sd39};
        weights3[6] = '{16'sd44, 16'sd108, 16'sd22, -16'sd225, 16'sd80, -16'sd194, 16'sd113, 16'sd59, 16'sd65, -16'sd259};
        weights3[7] = '{-16'sd64, 16'sd260, -16'sd138, -16'sd164, -16'sd100, 16'sd196, 16'sd223, -16'sd91, 16'sd79, 16'sd113};
        weights3[8] = '{16'sd81, -16'sd42, 16'sd89, -16'sd57, -16'sd207, -16'sd56, 16'sd26, -16'sd175, -16'sd16, -16'sd124};
        weights3[9] = '{-16'sd21, -16'sd270, -16'sd51, -16'sd167, 16'sd182, -16'sd186, 16'sd155, 16'sd96, 16'sd131, -16'sd6};
        weights3[10] = '{-16'sd167, 16'sd158, -16'sd130, 16'sd35, 16'sd142, 16'sd164, -16'sd34, -16'sd153, -16'sd20, -16'sd69};
        weights3[11] = '{16'sd90, 16'sd44, -16'sd10, -16'sd262, -16'sd100, 16'sd42, -16'sd228, -16'sd69, -16'sd19, 16'sd2};
        weights3[12] = '{-16'sd134, 16'sd31, 16'sd138, -16'sd92, -16'sd75, -16'sd221, -16'sd13, 16'sd117, -16'sd50, 16'sd115};
        weights3[13] = '{-16'sd241, 16'sd14, -16'sd15, -16'sd68, 16'sd205, -16'sd91, -16'sd59, 16'sd93, -16'sd294, 16'sd179};
        weights3[14] = '{-16'sd123, -16'sd175, 16'sd35, -16'sd127, -16'sd60, 16'sd70, -16'sd5, -16'sd215, 16'sd188, 16'sd96};
        weights3[15] = '{16'sd87, -16'sd62, 16'sd75, 16'sd183, -16'sd106, 16'sd159, 16'sd164, 16'sd10, -16'sd4, -16'sd156};
    end

    logic signed [15:0] layer1_out [N_LAYER1];
    logic signed [15:0] relu1_out [N_LAYER1];
    logic signed [15:0] layer2_out [N_LAYER2];
    logic signed [15:0] relu2_out [N_LAYER2];
    logic signed [15:0] layer3_out [N_LAYER3];

    // Layer 1: input -> matmul -> relu
    nn_layers #(.N_INPUTS(N_INPUTS), .N_OUTPUTS(N_LAYER1)) u_matmul1 (
        .input_vec(input_vec),
        .weights(weights1),
        .output_vec(layer1_out)
    );
    relu #(.N(N_LAYER1)) u_relu1 (
        .in_vec(layer1_out),
        .out_vec(relu1_out)
    );

    // Layer 2: relu1_out -> matmul -> relu
    nn_layers #(.N_INPUTS(N_LAYER1), .N_OUTPUTS(N_LAYER2)) u_matmul2 (
        .input_vec(relu1_out),
        .weights(weights2),
        .output_vec(layer2_out)
    );
    relu #(.N(N_LAYER2)) u_relu2 (
        .in_vec(layer2_out),
        .out_vec(relu2_out)
    );

    // Layer 3: relu2_out -> matmul -> argmax
    nn_layers #(.N_INPUTS(N_LAYER2), .N_OUTPUTS(N_LAYER3)) u_matmul3 (
        .input_vec(relu2_out),
        .weights(weights3),
        .output_vec(layer3_out)
    );
    argmax #(.N(N_LAYER3)) u_argmax (
        .in_vec(layer3_out),
        .pred(prediction)
    );
endmodule